`timescale 1ns/1ps

module system
(
  input wire CLK50MHZ,//GCLK
  /* input wire CLK32768KHZ,//RTC_CLK */

  input wire fpga_rst,//FPGA_RESET-T6
  input wire mcu_rst,//MCU_RESET-P20


  // Dedicated QSPI interface
  /*
  output wire qspi0_cs,
  output wire qspi0_sck,
  inout  wire [3:0] qspi0_dq,
  */
                           
  //gpioA
  // inout wire [31:0] gpioA,//GPIOA00~GPIOA31

  //gpioB
  // inout wire [31:0] gpioB,//GPIOB00~GPIOB31

  //uart0
  inout wire uart0_tx,
  inout wire uart0_rx,

  // JD (used for JTAG connection)
  inout wire mcu_TDO,//MCU_TDO-N17
  inout wire mcu_TCK,//MCU_TCK-P15 
  inout wire mcu_TDI,//MCU_TDI-T18
  inout wire mcu_TMS,//MCU_TMS-P17

  //pmu_wakeup(connected to LED)
  inout wire pmu_paden,  //PMU_VDDPADEN-U15
  inout wire pmu_padrst, //PMU_VADDPARST_V15
  inout wire mcu_wakeup  //MCU_WAKE-N15
);


  wire mmcm_locked;

  wire reset_periph;

  wire ck_rst;

  // All wires connected to the chip top
  wire dut_clock;
  wire dut_reset;

  wire dut_io_pads_jtag_TCK_i_ival;
  wire dut_io_pads_jtag_TMS_i_ival;
  wire dut_io_pads_jtag_TMS_o_oval;
  wire dut_io_pads_jtag_TMS_o_oe;
  wire dut_io_pads_jtag_TMS_o_ie;
  wire dut_io_pads_jtag_TMS_o_pue;
  wire dut_io_pads_jtag_TMS_o_ds;
  wire dut_io_pads_jtag_TDI_i_ival;
  wire dut_io_pads_jtag_TDO_o_oval;
  wire dut_io_pads_jtag_TDO_o_oe;

  wire [32-1:0] dut_io_pads_gpioA_i_ival;
  wire [32-1:0] dut_io_pads_gpioA_o_oval;
  wire [32-1:0] dut_io_pads_gpioA_o_oe;

  wire [32-1:0] dut_io_pads_gpioB_i_ival;
  wire [32-1:0] dut_io_pads_gpioB_o_oval;
  wire [32-1:0] dut_io_pads_gpioB_o_oe;

  wire dut_io_pads_qspi0_sck_o_oval;
  wire dut_io_pads_qspi0_cs_0_o_oval;
  wire dut_io_pads_qspi0_dq_0_i_ival;
  wire dut_io_pads_qspi0_dq_0_o_oval;
  wire dut_io_pads_qspi0_dq_0_o_oe;
  wire dut_io_pads_qspi0_dq_1_i_ival;
  wire dut_io_pads_qspi0_dq_1_o_oval;
  wire dut_io_pads_qspi0_dq_1_o_oe;
  wire dut_io_pads_qspi0_dq_2_i_ival;
  wire dut_io_pads_qspi0_dq_2_o_oval;
  wire dut_io_pads_qspi0_dq_2_o_oe;
  wire dut_io_pads_qspi0_dq_3_i_ival;
  wire dut_io_pads_qspi0_dq_3_o_oval;
  wire dut_io_pads_qspi0_dq_3_o_oe;


  wire dut_io_pads_aon_erst_n_i_ival;
  wire dut_io_pads_aon_pmu_dwakeup_n_i_ival;
  wire dut_io_pads_aon_pmu_vddpaden_o_oval;
  wire dut_io_pads_aon_pmu_padrst_o_oval ;
  wire dut_io_pads_bootrom_n_i_ival;
  wire dut_io_pads_dbgmode0_n_i_ival;
  wire dut_io_pads_dbgmode1_n_i_ival;
  wire dut_io_pads_dbgmode2_n_i_ival;

  //=================================================
  // Clock & Reset
  wire clk_16M;
  wire clk_8388608HZ;
  wire clk_32768HZ;


  mmcm ip_mmcm
  (
    .resetn(ck_rst),
    .clk_in(CLK50MHZ),
    
    .clk_out1(clk_16M),       // 16 MHz, this clock we set to core
    .clk_out2(clk_8388608HZ), // 32.768KHz, this clock we set to RTC

    .locked(mmcm_locked)
  );

  clk_div u_clk_div(
      .clk_in   ( clk_8388608HZ   ),
      .rst_n    ( ~ck_rst         ),
      .clk_out  ( clk_32768HZ     )
  );


  assign ck_rst = fpga_rst & mcu_rst;

  

  reset_sys ip_reset_sys
  (
    .slowest_sync_clk(clk_16M),
    .ext_reset_in(ck_rst), // Active-low
    .aux_reset_in(1'b1),
    .mb_debug_sys_rst(1'b0),
    .dcm_locked(mmcm_locked),
    .mb_reset(),
    .bus_struct_reset(),
    .peripheral_reset(reset_periph),
    .interconnect_aresetn(),
    .peripheral_aresetn()
  );


  //=================================================
  // UART0 Interface
 //* io_pads_gpioA_o_oval[16] <-> io_pads_uart0_rxd_o_oval;
 //* io_pads_gpioA_o_oval[17] <-> io_pads_uart0_txd_o_oval;
  wire       iobuf_uart0_rx_o;
  wire       iobuf_uart0_tx_o;

  IOBUF
  #(
    .DRIVE(12),             // Output drive strength set to 12 mA
    .IBUF_LOW_PWR("TRUE"),  // Enable low power mode for input buffer
    .IOSTANDARD("DEFAULT"), // Use default I/O standard
    .SLEW("SLOW")           // Set slew rate to slow for better signal integrity
  )
  iobuf_uart0_rx_o
  (
    .O(iobuf_uart0_rx_o),
    .IO(uart0_rx),                    // UART RX pin
    .I(dut_io_pads_gpioA_o_oval[16]), // No output from the FPGA
    .T(~dut_io_pads_gpioA_o_oe[16])   // Always drive high (input mode)
  );
  assign dut_io_pads_gpioA_i_ival[16] = iobuf_uart0_rx_o;

  IOBUF
  #(
    .DRIVE(12),             // Output drive strength set to 12 mA
    .IBUF_LOW_PWR("TRUE"),  // Enable low power mode for input buffer
    .IOSTANDARD("DEFAULT"), // Use default I/O standard
    .SLEW("SLOW")           // Set slew rate to slow for better signal integrity
  )
  iobuf_uart0_tx_o
  (
    .O(iobuf_uart0_tx_o),
    .IO(uart0_tx),                     // UART TX pin
    .I(dut_io_pads_gpioA_o_oval[17]),  // Output from the FPGA
    .T(~dut_io_pads_gpioA_o_oe[17])   // Drive low when output is enabled
  );


  //=================================================
  // SPI0 Interface
  // Declare wires for SPI0 data signals
  wire [3:0] qspi0_ui_dq_o;  // Output data from the e203 to the FPGA SPI Pins
  wire [3:0] qspi0_ui_dq_oe; // Output enable signals for SPI data lines
  wire [3:0] qspi0_ui_dq_i;  // Input data from the FPGA SPI Pins to the e203

  // Instantiate pull-up resistors for the SPI data lines
  // Ensures the lines are pulled to a high logic level when not driven
  // PULLUP qspi0_pullup[3:0]
  // (
  //   .O(qspi0_dq) // Connect to the bidirectional SPI data lines(qspi0_dq)
  // );

  // Instantiate IOBUFs for SPI data lines
  // IOBUFs allow bidirectional communication on the same physical pin
  // IOBUF qspi0_iobuf[3:0]
  // (
  //   .IO(qspi0_dq),        // Bidirectional SPI Pins
  //   .O(qspi0_ui_dq_i),    // Input data from FPGA SPI Pins to the e203
  //   .I(qspi0_ui_dq_o),    // Output data from e203 to FPGA SPI Pins
  //   .T(~qspi0_ui_dq_oe)   // High -> FPGA to e203, Low -> e203 to FPGA
  // );


  //=================================================
  // IOBUF instantiation for GPIOs
  /*
  IOBUF
  #(
    .DRIVE(12),             // Output drive strength set to 12 mA
    .IBUF_LOW_PWR("TRUE"),  // Enable low power mode for input buffer
    .IOSTANDARD("DEFAULT"), // Use default I/O standard
    .SLEW("SLOW")           // Set slew rate to slow for better signal integrity
  )
  gpioA_iobuf[31:0]
  (
    .O(dut_io_pads_gpioA_i_ival),
    .IO(gpioA),
    .I(dut_io_pads_gpioA_o_oval),
    .T(~dut_io_pads_gpioA_o_oe)
  );

  IOBUF
  #(
    .DRIVE(12),
    .IBUF_LOW_PWR("TRUE"),
    .IOSTANDARD("DEFAULT"),
    .SLEW("SLOW")
  )
  gpioB_iobuf[31:0]
  (
    .O(dut_io_pads_gpioB_i_ival),
    .IO(gpioB),
    .I(dut_io_pads_gpioB_o_oval),
    .T(~dut_io_pads_gpioB_o_oe)
  );
  */


  //=================================================
  // JTAG IOBUFs
  wire iobuf_jtag_TCK_o;
  IOBUF
  #(
    .DRIVE(12),
    .IBUF_LOW_PWR("TRUE"),
    .IOSTANDARD("DEFAULT"),
    .SLEW("SLOW")
  )
  IOBUF_jtag_TCK
  (
    .O(iobuf_jtag_TCK_o),
    .IO(mcu_TCK),
    .I(1'b0),
    .T(1'b1)
  );
  assign dut_io_pads_jtag_TCK_i_ival = iobuf_jtag_TCK_o ;
  PULLUP pullup_TCK (.O(mcu_TCK));

  wire iobuf_jtag_TMS_o;
  IOBUF
  #(
    .DRIVE(12),
    .IBUF_LOW_PWR("TRUE"),
    .IOSTANDARD("DEFAULT"),
    .SLEW("SLOW")
  )
  IOBUF_jtag_TMS
  (
    .O(iobuf_jtag_TMS_o),
    .IO(mcu_TMS),
    .I(1'b0),
    .T(1'b1)
  );
  assign dut_io_pads_jtag_TMS_i_ival = iobuf_jtag_TMS_o;
  PULLUP pullup_TMS (.O(mcu_TMS));

  wire iobuf_jtag_TDI_o;
  IOBUF
  #(
    .DRIVE(12),
    .IBUF_LOW_PWR("TRUE"),
    .IOSTANDARD("DEFAULT"),
    .SLEW("SLOW")
  )
  IOBUF_jtag_TDI
  (
    .O(iobuf_jtag_TDI_o),
    .IO(mcu_TDI),
    .I(1'b0),
    .T(1'b1)
  );
  assign dut_io_pads_jtag_TDI_i_ival = iobuf_jtag_TDI_o;
  PULLUP pullup_TDI (.O(mcu_TDI));

  wire iobuf_jtag_TDO_o;
  IOBUF
  #(
    .DRIVE(12),
    .IBUF_LOW_PWR("TRUE"),
    .IOSTANDARD("DEFAULT"),
    .SLEW("SLOW")
  )
  IOBUF_jtag_TDO
  (
    .O(iobuf_jtag_TDO_o),
    .IO(mcu_TDO),
    .I(dut_io_pads_jtag_TDO_o_oval),
    .T(~dut_io_pads_jtag_TDO_o_oe)
  );

  //! TRST is a optional pin for JTAG, not used in this design.
  //wire iobuf_jtag_TRST_n_o;
  //IOBUF
  //#(
  //  .DRIVE(12),
  //  .IBUF_LOW_PWR("TRUE"),
  //  .IOSTANDARD("DEFAULT"),
  //  .SLEW("SLOW")
  //)

  //=================================================
  // Assignment of IOBUF "IO" pins to package pins

  // Pins IO0-IO13
  // Shield header row 0: PD0-PD7

  // Use the LEDs for some more useful debugging things.
  assign pmu_paden  = dut_io_pads_aon_pmu_vddpaden_o_oval;  
  assign pmu_padrst = dut_io_pads_aon_pmu_padrst_o_oval;		

  // model select
  /*
  //* bootrom_n_i_ival: 0 = bootrom(0x0000_1000), 1 = flash(0x2000_0000)
  */
  assign dut_io_pads_bootrom_n_i_ival  = 1'b0;
  // assign dut_io_pads_bootrom_n_i_ival  = 1'b1;
  assign dut_io_pads_dbgmode0_n_i_ival = 1'b1;
  assign dut_io_pads_dbgmode1_n_i_ival = 1'b1;
  assign dut_io_pads_dbgmode2_n_i_ival = 1'b1;
  

  e203_soc_top dut
  (
    .hfextclk(clk_16M),
    .hfxoscen(),

    .lfextclk(clk_32768HZ), 
    .lfxoscen(),

    // Note: this is the real SoC top AON domain slow clock
    .io_pads_jtag_TCK_i_ival  (dut_io_pads_jtag_TCK_i_ival),
    .io_pads_jtag_TMS_i_ival  (dut_io_pads_jtag_TMS_i_ival),
    .io_pads_jtag_TDI_i_ival  (dut_io_pads_jtag_TDI_i_ival),
    .io_pads_jtag_TDO_o_oval  (dut_io_pads_jtag_TDO_o_oval),
    .io_pads_jtag_TDO_o_oe    (dut_io_pads_jtag_TDO_o_oe),

    .io_pads_gpioA_i_ival     (dut_io_pads_gpioA_i_ival),
    .io_pads_gpioA_o_oval     (dut_io_pads_gpioA_o_oval),
    .io_pads_gpioA_o_oe       (dut_io_pads_gpioA_o_oe),

    .io_pads_gpioB_i_ival     (dut_io_pads_gpioB_i_ival),
    .io_pads_gpioB_o_oval     (dut_io_pads_gpioB_o_oval),
    .io_pads_gpioB_o_oe       (dut_io_pads_gpioB_o_oe),

    .io_pads_qspi0_sck_o_oval (dut_io_pads_qspi0_sck_o_oval),
    .io_pads_qspi0_cs_0_o_oval(dut_io_pads_qspi0_cs_0_o_oval),

    .io_pads_qspi0_dq_0_i_ival(dut_io_pads_qspi0_dq_0_i_ival),
    .io_pads_qspi0_dq_0_o_oval(dut_io_pads_qspi0_dq_0_o_oval),
    .io_pads_qspi0_dq_0_o_oe  (dut_io_pads_qspi0_dq_0_o_oe),
    .io_pads_qspi0_dq_1_i_ival(dut_io_pads_qspi0_dq_1_i_ival),
    .io_pads_qspi0_dq_1_o_oval(dut_io_pads_qspi0_dq_1_o_oval),
    .io_pads_qspi0_dq_1_o_oe  (dut_io_pads_qspi0_dq_1_o_oe),
    .io_pads_qspi0_dq_2_i_ival(dut_io_pads_qspi0_dq_2_i_ival),
    .io_pads_qspi0_dq_2_o_oval(dut_io_pads_qspi0_dq_2_o_oval),
    .io_pads_qspi0_dq_2_o_oe  (dut_io_pads_qspi0_dq_2_o_oe),
    .io_pads_qspi0_dq_3_i_ival(dut_io_pads_qspi0_dq_3_i_ival),
    .io_pads_qspi0_dq_3_o_oval(dut_io_pads_qspi0_dq_3_o_oval),
    .io_pads_qspi0_dq_3_o_oe  (dut_io_pads_qspi0_dq_3_o_oe),


    //* Note: this is the real SoC top level reset signal
    .io_pads_aon_erst_n_i_ival       (ck_rst),
    .io_pads_aon_pmu_dwakeup_n_i_ival(dut_io_pads_aon_pmu_dwakeup_n_i_ival),
    .io_pads_aon_pmu_vddpaden_o_oval (dut_io_pads_aon_pmu_vddpaden_o_oval),
    .io_pads_aon_pmu_padrst_o_oval   (dut_io_pads_aon_pmu_padrst_o_oval ),

    .io_pads_bootrom_n_i_ival        (dut_io_pads_bootrom_n_i_ival),

    .io_pads_dbgmode0_n_i_ival       (dut_io_pads_dbgmode0_n_i_ival),
    .io_pads_dbgmode1_n_i_ival       (dut_io_pads_dbgmode1_n_i_ival),
    .io_pads_dbgmode2_n_i_ival       (dut_io_pads_dbgmode2_n_i_ival) 
  );

  // Assign reasonable values to otherwise unconnected inputs to chip top
  wire iobuf_dwakeup_o;
  IOBUF
  #(
    .DRIVE(12),
    .IBUF_LOW_PWR("TRUE"),
    .IOSTANDARD("DEFAULT"),
    .SLEW("SLOW")
  )
  IOBUF_dwakeup_n
  (
    .O(iobuf_dwakeup_o),
    .IO(mcu_wakeup),
    .I(1'b1),
    .T(1'b1)
  );
  assign dut_io_pads_aon_pmu_dwakeup_n_i_ival = (~iobuf_dwakeup_o);
  assign dut_io_pads_aon_pmu_vddpaden_i_ival  = 1'b1;

  /*
  assign qspi0_sck = dut_io_pads_qspi0_sck_o_oval;
  assign qspi0_cs  = dut_io_pads_qspi0_cs_0_o_oval;
  assign qspi0_ui_dq_o = {
    dut_io_pads_qspi0_dq_3_o_oval,
    dut_io_pads_qspi0_dq_2_o_oval,
    dut_io_pads_qspi0_dq_1_o_oval,
    dut_io_pads_qspi0_dq_0_o_oval
  };
  assign qspi0_ui_dq_oe = {
    dut_io_pads_qspi0_dq_3_o_oe,
    dut_io_pads_qspi0_dq_2_o_oe,
    dut_io_pads_qspi0_dq_1_o_oe,
    dut_io_pads_qspi0_dq_0_o_oe
  };
  assign dut_io_pads_qspi0_dq_0_i_ival = qspi0_ui_dq_i[0];
  assign dut_io_pads_qspi0_dq_1_i_ival = qspi0_ui_dq_i[1];
  assign dut_io_pads_qspi0_dq_2_i_ival = qspi0_ui_dq_i[2];
  assign dut_io_pads_qspi0_dq_3_i_ival = qspi0_ui_dq_i[3];
  */



endmodule


